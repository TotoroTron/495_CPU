library ieee;
use ieee.std_logic_1164.all;
library lpm;
use lpm.lpm_components.all;
use work.all;

entity cpu is
	port(
		clk : in std_logic
	);
end entity;

architecture dataflow of cpu is
begin
	

end architecture;