entity display is

end entity;

architecture behavioral of display is
begin


end architecture;