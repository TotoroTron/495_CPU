entity reg_file is
	port(
		clk : in std_logic;
	);
end entity;

architecture structural of reg_file is

begin


end architecture;